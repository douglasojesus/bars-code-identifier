library verilog;
use verilog.vl_types.all;
entity identificadorDeCodigoDeBarras_vlg_sample_tst is
    port(
        E0              : in     vl_logic;
        E1              : in     vl_logic;
        E2              : in     vl_logic;
        E3              : in     vl_logic;
        E4              : in     vl_logic;
        E5              : in     vl_logic;
        E6              : in     vl_logic;
        E7              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end identificadorDeCodigoDeBarras_vlg_sample_tst;

library verilog;
use verilog.vl_types.all;
entity identificadorDeCodigoDeBarras_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        L0              : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        L5              : in     vl_logic;
        L6              : in     vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        dig             : in     vl_logic;
        e               : in     vl_logic;
        f               : in     vl_logic;
        g               : in     vl_logic;
        ledG            : in     vl_logic;
        ledR            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end identificadorDeCodigoDeBarras_vlg_check_tst;
